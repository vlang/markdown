module native

fn to_html() string {
	return ''
}
