module native

struct Scanner {
}

fn new_scanner() Scanner {
	return Scanner{}
}
